* Selfmade model of the LM334 from National Semiconductor or ST
* Helmut Sennewald
*
* Pin order: v+  v-  R
.SUBCKT LM334 v+ v- R
Q4 N002 N001 v+ 0 pnp1
Q5 N003 N001 v+ 0 pnp1
Q6 R N001 v+ 0 pnp1 14
Q1 N003 N003 R 0 npn1 14
Q2 N002 N003 N004 0 npn1
Q3 N001 N002 R 0 npn1
C1 N002 N004 50p
R2 N004 v- 1ľ
R8 v+ v- 1G
C2 v+ v- 10p
C3 N003 v- 1p
C4 R v- 1p
.model npn1 NPN(Is=1e-15 BF=200 TF=1e-9 Cjc=0.5e-12 Cje=1e-12 VAF=100 Rb=100 Re=5)
.model pnp1 PNP(Is=1e-15 BF=100 TF=1e-7 Cjc=0.5e-12 Cje=1e-12 VAF=100 Rb=100 Re=5)
.ENDS